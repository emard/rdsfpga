../fmgen.vhd