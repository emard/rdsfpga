--
-- Copyright (c) 2013 - 2015 Marko Zec, University of Zagreb
-- Copyright (c) 2015 Davor Jadrijevic
-- All rights reserved.
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in the
--    documentation and/or other materials provided with the distribution.
--
-- THIS SOFTWARE IS PROVIDED BY THE AUTHOR AND CONTRIBUTORS ``AS IS'' AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
-- ARE DISCLAIMED.  IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE LIABLE
-- FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
-- DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
-- LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
-- OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
-- SUCH DAMAGE.
--
-- $Id$
--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

use work.message.all; -- RDS message in file message.vhd

entity bram_rds is
    port(
	clk: in std_logic;
	imem_addr: in std_logic_vector(8 downto 0);
	imem_data_out: out std_logic_vector(7 downto 0)
--	dmem_write: in std_logic;
--	dmem_byte_sel: in std_logic_vector(3 downto 0);
--	dmem_addr: in std_logic_vector(31 downto 2);
--	dmem_data_in: in std_logic_vector(7 downto 0);
--	dmem_data_out: out std_logic_vector(7 downto 0)
    );
end bram_rds;

architecture x of bram_rds is
   signal bram_0: rds_msg_type := rds_msg_map;
   signal ibram_0: std_logic_vector(7 downto 0);
begin
   imem_data_out <= ibram_0;

--   process(clk)
--   begin
--	if falling_edge(clk) then
--	  ibram_0 <= bram_0(conv_integer(imem_addr));
--	end if;
--   end process;

   ibram_0 <= bram_0(conv_integer(imem_addr));
end x;
