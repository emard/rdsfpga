message-hello.vhd