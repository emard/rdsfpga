../lattice/lattice_pll_25MHz_250MHz.vhd