../enkoder.vhd