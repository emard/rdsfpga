../tonegen-rds.vhd