message-custom.vhd